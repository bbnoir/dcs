../01_RTL/Seq.sv