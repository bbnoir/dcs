../00_TESTBED/testbench1.sv