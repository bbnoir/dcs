../01_RTL/DCT.sv