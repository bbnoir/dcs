../01_RTL/HE.sv