../00_TESTBED/testbench5.sv