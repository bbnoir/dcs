../01_RTL/Counter.sv