../01_RTL/CDC.sv