../01_RTL/Sort.sv