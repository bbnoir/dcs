../00_TESTBED/pattern.sv