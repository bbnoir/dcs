../01_RTL/TL.sv