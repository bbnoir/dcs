../01_RTL/SMJ.sv