/RAID2/COURSE/dcs/dcs064/Lab02/01_RTL/Bubble.sv