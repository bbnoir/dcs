../00_TESTBED/testbench4.sv