/RAID2/COURSE/dcs/dcs064/Lab06/00_TESTBED/pattern.sv