../01_RTL/P_MUL.sv