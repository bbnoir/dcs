../01_RTL/mem_slave.sv