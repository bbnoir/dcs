../00_TESTBED/testbench3.sv