../00_TESTBED/testbench2.sv