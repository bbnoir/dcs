../00_TESTBED/testbench.sv