../01_RTL/MIPS.sv