../00_TESTBED/testbench6.sv