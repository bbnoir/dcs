../01_RTL/inter.sv