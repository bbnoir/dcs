../01_RTL/Fpc.sv