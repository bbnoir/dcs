../00_TESTBED/TESTBENCH.sv