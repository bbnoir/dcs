../02_SYN/Netlist/SS_SYN.sv