../01_RTL/I2S.sv