../01_RTL/BCD.sv